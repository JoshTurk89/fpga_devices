
------------------------------------------------------------------------------
-- Device/Project:  Testbench Device/Project name
-- File: 	          tb_dev_prj.vhd
-- Author:	        Joshua Jesus Quintana Di­az
-- Date:	          dd/mm/yy
-- Version:	        1.0
-- History:	        1.0 Initial Version
------------------------------------------------------------------------------
-- Description: 
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.log2;
use ieee.math_real.ceil;
use ieee.math_real.floor;

library work;
use work.logger_pkg.all;
use work.tb_common_pkg.all;
use work.test000000.all;

entity tb_device_project_arch is
  generic (g_numtest : string(1 to 6) := "000000"
                                         );
end tb_device_project_arch;

architecture beh of tb_device_project_arch is

  -----------------------------------------------------------------------------------------
  -- --------------------------- TEST CLKS SIGNALS ----------------------------------------
  -----------------------------------------------------------------------------------------
  signal tb_clk             : std_logic := '1';
  signal tb_reset_n         : std_logic;

  --------------------------------------------------------------------------------
  --------------------- CONSTANT -------------------------------------------------
  --------------------------------------------------------------------------------

  --------------------------------------------------------------------------------
  ---------------------- TYPES ---------------------------------------------------
  --------------------------------------------------------------------------------

  --------------------------------------------------------------------------------
  ------------------- TEST SIGNALS -----------------------------------------------
  --------------------------------------------------------------------------------

  --------------------------------------------------------------------------------
  -------------- SEQUENCES SIGNALS -----------------------------------------------
  --------------------------------------------------------------------------------
  signal tb_sq_start        : std_logic;
  signal tb_sq_busy         : std_logic;

begin

  p_stimuli : process
  begin
    case g_numtest is
      when "000000" => test000000_example (tb_clk, tb_reset_n, tb_sq_start, tb_sq_busy);
      when others => assert false report "test " & g_numtest & " not defined" severity failure;
    end case;
    wait;
  end process p_stimuli;

  -------------------------------------------------------------------------------- 
  ------------------------ Clk generations ---------------------------------------
  --------------------------------------------------------------------------------
  tb_clk     <= not(tb_clk) after C_CLK_SYS/2;

  --------------------------------------------------------------------------------
  ------------------------ rst generations ---------------------------------------
  --------------------------------------------------------------------------------
  tb_reset_n <= '0', '1' after 200 ns;

  --------------------------------------------------------------------------------
  ------------------ DUT COMPONENT INSTANTIATION ---------------------------------
  --------------------------------------------------------------------------------  

  DUT : device
  generic map(
    G_example_1 => example_1,
    G_example_2 => example_2
  )
  port map(
    EXAMPLE_1 => example_1,
    EXAMPLE_2 => example_2
  );

  --------------------------------------------------------------------------------
  ----------------- AGENT COMPONENT INSTANTIATION --------------------------------
  -------------------------------------------------------------------------------- 
  ag_dev : device
  generic map(
    G_example_1 => example_1,
    G_example_2 => example_2
  )
  port map(
    EXAMPLE_1 => example_1,
    EXAMPLE_2 => example_2
  );

end beh;