
------------------------------------------------------------------------------
-- Device/Project: Logic Adder Device
-- File: 	device_project_arch_pkg.vhd
-- Author:	Joshua Jesus Quintana Di­az
-- Date:	
-- Version:	1.0
-- History:	1.0 Initial Version
-- Design:	
------------------------------------------------------------------------------
-- Description: 
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.log2;
use ieee.math_real.ceil;
use ieee.math_real.floor;

library work;
use work.TBD.all;

package device_project_arch_pkg is

  --------------------------------------------------------------------------------
  ---------------------- CONSTANT ------------------------------------------------
  --------------------------------------------------------------------------------

  --------------------------------------------------------------------------------
  ---------------------- TYPES ---------------------------------------------------
  --------------------------------------------------------------------------------

  --------------------------------------------------------------------------------
  ---------------------- PROCEDURES ----------------------------------------------
  --------------------------------------------------------------------------------
  procedure name_proc (
    constant C_1    : in  natural;
    constant C_2    : in  natural;
    variable v_1    : in  integer;
    variable v_2    : out integer;
    signal SIGNAL_1 : in  std_logic;
    signal SIGNAL_2 : out std_logic
  );

  --------------------------------------------------------------------------------
  ---------------------- FUNCTIONS -----------------------------------------------
  --------------------------------------------------------------------------------
  function name_func(entry_1 : integer; entry_2 : integer; entry_3 : std_logic) return std_logic_vector;

  --------------------------------------------------------------------------------
  ---------------------- COMPONENTS ----------------------------------------------
  --------------------------------------------------------------------------------  

  component device_project_arch is
    generic (

    );
    port (

    );
  end component;

end device_project_arch_pkg;

package body device_project_arch_pkg is

  --------------------------------------------------------------------------------
  ---------------------- PROCEDURES ----------------------------------------------
  --------------------------------------------------------------------------------
  procedure name_proc (
    constant C_1    : in  natural;
    constant C_2    : in  natural;
    variable v_1    : in  integer;
    variable v_2    : out integer;
    signal SIGNAL_1 : in  std_logic;
    signal SIGNAL_2 : out std_logic
  ) is    
  begin

    --------------------------------------------------------------------------------
    --------------------- I/O PROCEDURES -------------------------------------------
    --------------------------------------------------------------------------------

    --------------------------------------------------------------------------------
    --------------------- BODY -----------------------------------------------------
    --------------------------------------------------------------------------------

  end name_proc;

  --------------------------------------------------------------------------------
  ---------------------- FUNCTIONS -----------------------------------------------
  --------------------------------------------------------------------------------
  function name_func(entry_1 : integer; entry_2 : integer; entry_3 : std_logic) return std_logic_vector is
    variable v_example1 : std_logic_vector(entry_2 - 1 downto 0) := (others => '0');
  begin

    return std_logic_vector;

  end function;

end device_project_arch_pkg;
